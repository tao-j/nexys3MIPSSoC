`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:46:42 07/01/2012 
// Design Name: 
// Module Name:    Device_7seg 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module seven_seg_Dev_IO( input clk,
							input rst,
							input GPIOe0000000_we,
							input [2:0] Test,
							input [31:0] disp_cpudata,
							input [31:0] Test_data0,
							input [31:0] Test_data1,
							input [31:0] Test_data2,
							input [31:0] Test_data3,
							input [31:0] Test_data4,
							input [31:0] Test_data5,
							input [31:0] Test_data6,						 						 
							output[31:0] disp_num						 
						);

endmodule
